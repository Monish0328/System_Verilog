task (input sum[7:0] a,b output [7:0]c);
  begin 
    c=a+b;
  end
endtask
